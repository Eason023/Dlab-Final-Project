// physic.v
//-----------------------------------------------------------------------------
// �Ҳե\��G�M�`��֥d�C���Ʋy�C�������i�y�骫�z�B�ʡj�M�i�o���P�w�j�C
// �B�z�y����m�B�t�סB���O�B���ҸI���M����I���᪺�ϼu�p��C
// �ѪR�ץؼСG320 x 240
//-----------------------------------------------------------------------------

module physic (
    input wire clk,
    input wire rst_n,

    // P1 & P2 �ʧ@��J (�ȱ����ާ@�A�Ω����y�P�_)
    input wire p1_op_move_left, input wire p1_op_move_right, input wire p1_op_jump,
    input wire p2_op_move_left, input wire p2_op_move_right, input wire p2_op_jump,

    // �I���������G��J (�Ӧ� render/bounding detect �Ҳ�)
    input wire p1_cover, // P1 ���a�P�y�O�_�o�͸I��
    input wire p2_cover, // P2 ���a�P�y�O�_�o�͸I��
    
    // ���a����e��m (�ȥΩ�p�����y�᪺�y��_�l��m)
    // �O�� [9:0] ��e�A���ȷ|����b 0-320/240 �d��
    input wire [9:0] p1_pos_x_i, p1_pos_y_i,
    input wire [9:0] p2_pos_x_i, p2_pos_y_i,

    //-----------------------------------------------------
    // Output: ��X�y����e��m�M�C�����A
    //-----------------------------------------------------
    output reg [9:0] ball_pos_x, ball_pos_y,
    
    output reg [3:0] p1_score, p2_score,
    output reg game_over // �C���O�_���� (���o��/�y���a)
);
    
    //��e�w�q
    localparam COORD_W = 10; // �y�Ц�e (0-1023), ��ڨϥ� 0-320/240
    localparam VEL_W   = 10; // �t�צ�e (�w�I�� Q4.6)
    localparam FRAC_W  = 6;  // �w�I�ƪ��p�Ƴ�����e
    localparam SCORE_W = 4;  // ���Ʀ�e (0-15)

    //���z�`�� (�w�I�� Q4.6: 1.0 = 10'd64)
    localparam FRAC_ONE = 10'd64; 
    localparam GRAVITY = 10'd2;   
    localparam BOUNCE_DAMPING = 10'd55; 

    //���y�ϼu�t��
    localparam P1_HIT_VX = 10'd192; 
    localparam P1_HIT_VY = 10'd320; 
    localparam P2_HIT_VX = -10'd192; 
    localparam P2_HIT_VY = 10'd320; 

    localparam SCREEN_WIDTH = 10'd320;
    localparam SCREEN_HEIGHT = 10'd240;

    localparam NET_X_POS = 10'd160;     // �y�� X �y�� (���u 320/2)
    localparam NET_W = 10'd6;           // �y���b�e (�z�n�D���Ѽ�)
    localparam NET_H = 10'd90;          // �y������ (�z�n�D���Ѽ�)
    localparam FLOOR_Y_POS = 10'd30;    // �a�� Y �y�� (�۹���C)
    
    localparam NET_TOP_Y = FLOOR_Y_POS + NET_H; // �y������ Y �y��

    localparam LEFT_WALL_X = 10'd0;
    localparam RIGHT_WALL_X = SCREEN_WIDTH - 1; // 319

    localparam BALL_INIT_X = NET_X_POS;
    localparam BALL_INIT_Y = 10'd150; // �e�����u���W
    
    reg [VEL_W-1:0] ball_vel_x, ball_vel_y;
    
    wire [VEL_W-1:0] ball_vel_y_calc; 
    wire [COORD_W-1:0] ball_pos_y_calc;
    
    wire ball_hit_floor_p1_side; 
    wire ball_hit_floor_p2_side; 
    
    // �s�W���l�����I��
    wire ball_hit_net_top;
    // �ק���l�����I��
    wire ball_hit_net_side_p1;
    wire ball_hit_net_side_p2;

    wire ball_hit_wall_side;     
    
    //1. ���z�B�ʾǭp�� (�U�@�g���w�p���A)

    assign ball_vel_y_calc = ball_vel_y - GRAVITY; 
    assign ball_pos_y_calc = ball_pos_y + (ball_vel_y_calc >>> FRAC_W);
    
    //2. ���ҸI���P�o������

    // �y���a/�o������ (�y�� Y �y�Фp�󵥩�a�� Y �y��)
    assign ball_hit_floor_p1_side = (ball_pos_y_calc <= FLOOR_Y_POS) && (ball_pos_x_calc < NET_X_POS);
    assign ball_hit_floor_p2_side = (ball_pos_y_calc <= FLOOR_Y_POS) && (ball_pos_x_calc >= NET_X_POS);

    // ���lX�b�d��P�_
    wire ball_in_net_x_range = (ball_pos_x < NET_X_POS + NET_W) && (ball_pos_x > NET_X_POS - NET_W);

    // ���l�����I�� (�q�W��{�����)
    assign ball_hit_net_top = ball_in_net_x_range && 
                              (ball_pos_y > NET_TOP_Y) &&           // ��e�b�����W��
                              (ball_pos_y_calc <= NET_TOP_Y);       // �U�@�g���������

    // ���l�����I�� (������l�D��A�ư�����)
    assign ball_hit_net_side_p1 = ball_in_net_x_range && 
                                  (ball_pos_x_calc < NET_X_POS) &&  // �y�ߦb P1 ��
                                  (ball_pos_y_calc <= NET_TOP_Y) && // �B���צb���l�D�餺
                                  (ball_pos_y_calc > FLOOR_Y_POS);

    assign ball_hit_net_side_p2 = ball_in_net_x_range && 
                                  (ball_pos_x_calc >= NET_X_POS) && // �y�ߦb P2 ��
                                  (ball_pos_y_calc <= NET_TOP_Y) && // �B���צb���l�D�餺
                                  (ball_pos_y_calc > FLOOR_Y_POS);
                                  
    // ����I��
    assign ball_hit_wall_side = (ball_pos_x_calc <= LEFT_WALL_X) || (ball_pos_x_calc >= RIGHT_WALL_X);
    
    //3. �I�������P���A��s (�֤߲զX�޿�)
    
    reg [VEL_W-1:0] final_vel_x, final_vel_y;
    reg [COORD_W-1:0] final_pos_x, final_pos_y;
    reg [SCORE_W-1:0] p1_score_next, p2_score_next;
    
    reg score_happened; 
    
    assign game_over = score_happened; 

    always @(*) begin
        // �w�]�U�@���A
        final_vel_x = ball_vel_x;
        final_vel_y = ball_vel_y_calc;
        final_pos_x = ball_pos_x + (ball_vel_x >>> FRAC_W);
        final_pos_y = ball_pos_y_calc;
        
        p1_score_next = p1_score;
        p2_score_next = p2_score;
        score_happened = 1'b0; 

        // A. �u���ų̰����I���G�������y (�~����J p1_cover/p2_cover)
        if (p1_cover || p2_cover) begin
            if (p1_cover) begin
                final_vel_x = P1_HIT_VX;
                final_vel_y = P1_HIT_VY;
                final_pos_x = p1_pos_x_i + 30; // �T�O���d�I
                final_pos_y = p1_pos_y_i + 30;
            end
            else if (p2_cover) begin
                final_vel_x = P2_HIT_VX;
                final_vel_y = P2_HIT_VY;
                final_pos_x = p2_pos_x_i - 30; // �T�O���d�I
                final_pos_y = p2_pos_y_i + 30;
            end
        end
        // B. ���һP�o���I�� (�����B�z)
        else begin
            // 1. �o�����a (�̰��u���Ū����ҸI��)
            if (ball_hit_floor_p1_side) begin // �y���b P1 �ϡAP2 �o��
                p2_score_next = p2_score + 1;
                score_happened = 1'b1; 
            end 
            else if (ball_hit_floor_p2_side) begin // �y���b P2 �ϡAP1 �o��
                p1_score_next = p1_score + 1;
                score_happened = 1'b1; 
            end
            
            // 2. ���l�����I�� (�q�W�踨����l�W)
            else if (ball_hit_net_top) begin
                final_vel_y = (~final_vel_y + 1); // �����t�פϦV
                final_pos_y = NET_TOP_Y;         // ��w�b����
            end

            // 3. ���l�����I��
            else if (ball_hit_net_side_p1 || ball_hit_net_side_p2) begin
                final_vel_x = (~final_vel_x + 1); // �����t�פϦV
                // ��w��m�H�����z
                if (ball_pos_x_calc < NET_X_POS) final_pos_x = NET_X_POS - NET_W; // P1 ���ϼu
                else final_pos_x = NET_X_POS + NET_W;                           // P2 ���ϼu
            end

            // 4. �a���I�� (�D�o���ϡA�Y�Ʋy���U)
            else if (ball_pos_y_calc <= FLOOR_Y_POS) begin
                // �t�פϦV * �I��
                final_vel_y = (FRAC_ONE - ball_vel_y_calc) * BOUNCE_DAMPING / FRAC_ONE;
                final_pos_y = FLOOR_Y_POS; 
            end

            // 5. ����I��
            else if (ball_hit_wall_side) begin
                final_vel_x = (~final_vel_x + 1); 
                if (ball_pos_x_calc <= LEFT_WALL_X) final_pos_x = LEFT_WALL_X;
                if (ball_pos_x_calc >= RIGHT_WALL_X) final_pos_x = RIGHT_WALL_X;
            end
        end
    end

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            // �t�έ��m (�w�魫�m/�C�����})
            ball_pos_x <= BALL_INIT_X; ball_pos_y <= BALL_INIT_Y;
            ball_vel_x <= 0; ball_vel_y <= 0;
            p1_score <= 0; p2_score <= 0;
        end else begin
            
            // ���Ƨ�s
            p1_score <= p1_score_next;
            p2_score <= p2_score_next;

            //�y����m�M�t�ק�s (�p�G�o���A�h���m�y)
            if (score_happened) begin
                // �y�o��/�o�y���m�ɪ���m/�t��
                ball_pos_x <= BALL_INIT_X; 
                ball_pos_y <= BALL_INIT_Y;
                ball_vel_x <= 0;
                ball_vel_y <= 0;
            end else begin
                // ���`���z�B��
                ball_vel_x <= final_vel_x;
                ball_vel_y <= final_vel_y;
                ball_pos_x <= final_pos_x;
                ball_pos_y <= final_pos_y;
            end
        end
    end
endmodule